//
module pwm_core_ip();

endmodule