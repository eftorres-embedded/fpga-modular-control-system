module pwm_compare()

endmodule