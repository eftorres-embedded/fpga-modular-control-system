//uart_rx_engine.sv

module uart_rx_engine()







endmodule