module pwm_timebase()


endmodule